module Adder(input [31:0] in, pluser, output [31:0] out);
    assign out = in + pluser;
endmodule